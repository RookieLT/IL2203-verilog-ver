library verilog;
use verilog.vl_types.all;
entity tb_alu1 is
end tb_alu1;
