`timescale 1ns/1ns
module tb_microcontroller;

reg clk,rst;
reg [15:0] din;
wire rw;
wire [15:0] addr;
wire [15:0] dout;

microcontroller#(3,16) mc(din,clk,rst,rw,addr,dout);

initial clk=0;
always #2 clk=~clk;

initial begin
    rst<=1;
    // #10 rst <= 0;
    //     din <= 16'b1010_001_000000010;          //LDI
    // #20 din <= 16'b1010_101_100000000;          //LDI
    // #20 din <= 16'b1010_000_000000010;
    // //ADD
    // #20 din <= 16'b0000_011_101_001_000;
    // //SUB
    // #20 din <= 16'b0001_011_000_001_000;
    // //AND
    // #20 din <= 16'b0010_011_000_101_000;
    // //OR
    // #20 din <= 16'b0011_011_101_001_000;
    // //XOR
    // #20 din <= 16'b0100_011_101_001_000;
    // //NOT
    // #20 din <= 16'b0101_011_001_000_000;
    // //MOV
    // #20 din <= 16'b0110_011_101_000_000;
    // //NOP
    // #20 din <= 16'b0111_000_000_000_000;
    // //LD
    // #20 din <= 16'b1000_011_001_000_000;
    // #8 din <= 16'b0000_1111_0000_1111;
    // //ST
    // #12 din <= 16'b1001_000_001_101_000;
    // //NU
    // #20 din <= 16'b1011_000_000_000_000;
    // //BRZ
    // #20 din <= 16'b0001_011_000_001_000;
    // #20 din <= 16'b1100_000_000_111_111;
    // //BRN
    // #20 din <= 16'b0001_011_101_001_000;
    // #20 din <= 16'b1101_000_001_000_000;
    // //BRO
    // #20 din <= 16'b1010_010_100000000;
    // #20 din <= 16'b1110_000_000_111;
    // //BRA
    // #20 din <= 16'b1111_000_110_000_000;
    // #20 din <= 'b0;
end

endmodule